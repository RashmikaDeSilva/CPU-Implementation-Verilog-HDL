`timescale 1ns/100ps

// 2 to 1 multiplexer needed for Barrel Shifter
module MUX_2x1 (INPUT1, INPUT2, OUTPUT, SELECT );
    input INPUT1, INPUT2, SELECT;
    output wire OUTPUT;

    assign OUTPUT = (SELECT) ? INPUT1 : INPUT2;
endmodule

// Barrel shifter module for logical left shift
module barrelShifter_LSL( INPUT, SHIFTED_OUTPUT, SHIFT_AMOUNT);        

  input  [7:0] INPUT;                   //The 8-bit Input line 
  output  [7:0] SHIFTED_OUTPUT;         //The 8-bit Output line 
  input [2:0] SHIFT_AMOUNT;             //The 3-bit shift distance selection Input 
  wire [7:0] INTERIM_1,INTERIM_2;       //Two 8-bit intermediate lines 

  //the barrel shifter implemented as array of MUX s in 3 columns and 8 rows

  // MUX naming convetion :- MUX_CiRi - 2x1 MUX in i'th column and i'th row ; i = 0,1,2,3,4,5,6,7

  MUX_2x1 MUX_C0R0 (1'b0,  INPUT[0], INTERIM_1[0], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R1 (INPUT[0], INPUT[1], INTERIM_1[1], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R2 (INPUT[1], INPUT[2], INTERIM_1[2], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R3 (INPUT[2], INPUT[3], INTERIM_1[3], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R4 (INPUT[3], INPUT[4], INTERIM_1[4], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R5 (INPUT[4], INPUT[5], INTERIM_1[5], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R6 (INPUT[5], INPUT[6], INTERIM_1[6], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R7 (INPUT[6], INPUT[7], INTERIM_1[7], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C1R0 (1'b0  , INTERIM_1[0], INTERIM_2[0], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R1 (1'b0  , INTERIM_1[1], INTERIM_2[1], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R2 (INTERIM_1[0], INTERIM_1[2], INTERIM_2[2], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R3 (INTERIM_1[1], INTERIM_1[3], INTERIM_2[3], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R4 (INTERIM_1[2], INTERIM_1[4], INTERIM_2[4], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R5 (INTERIM_1[3], INTERIM_1[5], INTERIM_2[5], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R6 (INTERIM_1[4], INTERIM_1[6], INTERIM_2[6], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R7 (INTERIM_1[5], INTERIM_1[7], INTERIM_2[7], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C2R0 (1'b0  , INTERIM_2[0], SHIFTED_OUTPUT[0], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R1 (1'b0  , INTERIM_2[1], SHIFTED_OUTPUT[1], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R2 (1'b0  , INTERIM_2[2], SHIFTED_OUTPUT[2], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R3 (1'b0  , INTERIM_2[3], SHIFTED_OUTPUT[3], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R4 (INTERIM_2[0], INTERIM_2[4], SHIFTED_OUTPUT[4], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R5 (INTERIM_2[1], INTERIM_2[5], SHIFTED_OUTPUT[5], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R6 (INTERIM_2[2], INTERIM_2[6], SHIFTED_OUTPUT[6], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R7 (INTERIM_2[3], INTERIM_2[7], SHIFTED_OUTPUT[7], SHIFT_AMOUNT[2]); 

endmodule


// Barrel shifter module for logical right shift
module barrelShifter_LSR( INPUT, SHIFTED_OUTPUT, SHIFT_AMOUNT);        

  input  [7:0] INPUT;                   //The 8-bit Input line 
  output  [7:0] SHIFTED_OUTPUT;         //The 8-bit Output line 
  input [2:0] SHIFT_AMOUNT;             //The 3-bit shift magnitude selection Input 
  wire [7:0] INTERIM_1,INTERIM_2;       //Two 8-bit intermediate lines 

  //the barrel shifter implemented as array of MUX s in 3 columns and 8 rows

  // MUX naming convetion :- MUX_CiRi - 2x1 MUX in i'th column and i'th row ; i = 0,1,2,3,4,5,6,7 
  
  MUX_2x1 MUX_C0R0 (1'b0,  INPUT[7], INTERIM_1[0], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R1 (INPUT[7], INPUT[6], INTERIM_1[1], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R2 (INPUT[6], INPUT[5], INTERIM_1[2], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R3 (INPUT[5], INPUT[4], INTERIM_1[3], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R4 (INPUT[4], INPUT[3], INTERIM_1[4], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R5 (INPUT[3], INPUT[2], INTERIM_1[5], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R6 (INPUT[2], INPUT[1], INTERIM_1[6], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R7 (INPUT[1], INPUT[0], INTERIM_1[7], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C1R0 (1'b0  , INTERIM_1[0], INTERIM_2[0], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R1 (1'b0  , INTERIM_1[1], INTERIM_2[1], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R2 (INTERIM_1[0], INTERIM_1[2], INTERIM_2[2], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R3 (INTERIM_1[1], INTERIM_1[3], INTERIM_2[3], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R4 (INTERIM_1[2], INTERIM_1[4], INTERIM_2[4], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R5 (INTERIM_1[3], INTERIM_1[5], INTERIM_2[5], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R6 (INTERIM_1[4], INTERIM_1[6], INTERIM_2[6], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R7 (INTERIM_1[5], INTERIM_1[7], INTERIM_2[7], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C2R0 (1'b0  , INTERIM_2[0], SHIFTED_OUTPUT[7], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R1 (1'b0  , INTERIM_2[1], SHIFTED_OUTPUT[6], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R2 (1'b0  , INTERIM_2[2], SHIFTED_OUTPUT[5], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R3 (1'b0  , INTERIM_2[3], SHIFTED_OUTPUT[4], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R4 (INTERIM_2[0], INTERIM_2[4], SHIFTED_OUTPUT[3], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R5 (INTERIM_2[1], INTERIM_2[5], SHIFTED_OUTPUT[2], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R6 (INTERIM_2[2], INTERIM_2[6], SHIFTED_OUTPUT[1], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R7 (INTERIM_2[3], INTERIM_2[7], SHIFTED_OUTPUT[0], SHIFT_AMOUNT[2]); 

endmodule


// Barrel shifter module for arithmetic right shift
module barrelShifter_ASR( INPUT, SHIFTED_OUTPUT, SHIFT_AMOUNT);        

  input  [7:0] INPUT;                   //The 8-bit Input line 
  output  [7:0] SHIFTED_OUTPUT;         //The 8-bit Output line 
  input [2:0] SHIFT_AMOUNT;             //The 3-bit shift magnitude selection Input 
  wire [7:0] INTERIM_1,INTERIM_2;       //Two 8-bit intermediate lines 

  //the barrel shifter implemented as array of MUX s in 3 columns and 8 rows

  // MUX naming convetion :- MUX_CiRi - 2x1 MUX in i'th column and i'th row ; i = 0,1,2,3,4,5,6,7
  
  MUX_2x1 MUX_C0R0 (INPUT[7],  INPUT[7], INTERIM_1[0], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R1 (INPUT[7], INPUT[6], INTERIM_1[1], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R2 (INPUT[6], INPUT[5], INTERIM_1[2], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R3 (INPUT[5], INPUT[4], INTERIM_1[3], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R4 (INPUT[4], INPUT[3], INTERIM_1[4], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R5 (INPUT[3], INPUT[2], INTERIM_1[5], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R6 (INPUT[2], INPUT[1], INTERIM_1[6], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C0R7 (INPUT[1], INPUT[0], INTERIM_1[7], SHIFT_AMOUNT[0]); 

  MUX_2x1 MUX_C1R0 (INPUT[7], INTERIM_1[0], INTERIM_2[0], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R1 (INPUT[7], INTERIM_1[1], INTERIM_2[1], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R2 (INTERIM_1[0], INTERIM_1[2], INTERIM_2[2], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R3 (INTERIM_1[1], INTERIM_1[3], INTERIM_2[3], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R4 (INTERIM_1[2], INTERIM_1[4], INTERIM_2[4], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R5 (INTERIM_1[3], INTERIM_1[5], INTERIM_2[5], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R6 (INTERIM_1[4], INTERIM_1[6], INTERIM_2[6], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C1R7 (INTERIM_1[5], INTERIM_1[7], INTERIM_2[7], SHIFT_AMOUNT[1]); 

  MUX_2x1 MUX_C2R0 (INPUT[7], INTERIM_2[0], SHIFTED_OUTPUT[7], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R1 (INPUT[7], INTERIM_2[1], SHIFTED_OUTPUT[6], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R2 (INPUT[7], INTERIM_2[2], SHIFTED_OUTPUT[5], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R3 (INPUT[7], INTERIM_2[3], SHIFTED_OUTPUT[4], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R4 (INTERIM_2[0], INTERIM_2[4], SHIFTED_OUTPUT[3], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R5 (INTERIM_2[1], INTERIM_2[5], SHIFTED_OUTPUT[2], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R6 (INTERIM_2[2], INTERIM_2[6], SHIFTED_OUTPUT[1], SHIFT_AMOUNT[2]); 

  MUX_2x1 MUX_C2R7 (INTERIM_2[3], INTERIM_2[7], SHIFTED_OUTPUT[0], SHIFT_AMOUNT[2]); 

endmodule